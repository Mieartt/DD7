library ieee;
use ieee.std_logic_1164.all;
entity salah is
 port (
        fom    : in std_logic;
        khcham : out std_logic
 );
 end entity;
 architecture arch of salah is 
 begin
 end behavior;

 